module dmac_channel_requester (
    input clk,
    input rst
);

endmodule : dmac_channel_requester